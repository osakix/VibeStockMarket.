module vibe;
initial begin
  $display("Welcome to VibeStockMarket!");
  $finish;
end
endmodule
