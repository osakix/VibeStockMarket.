library ieee;
use ieee.std_logic_1164.all;
entity vibe is
end entity;
architecture behav of vibe is
begin
    process begin
        report "Welcome to VibeStockMarket!";
        wait;
    end process;
end architecture;
